package alu_pkg;
    import uvm_pkg ::*;
    `include "uvm_macros.svh"
    `include "sequence_item.svh"
     typedef uvm_sequencer#(sequence_item) sequencer;
    
    `include "result_transaction.svh"
    `include "scoreboard.svh"
    `include "command_monitor.svh"
    `include "result_monitor.svh"
    `include "driver.svh"
    `include "config_agent.svh"
    `include "agent.svh"
    `include "env.svh"    
    `include "base_test.svh"
    `include "reset_sequence.svh"
    `include "mode_a_sequence.svh"
    `include "mode_b_sequence.svh"
    `include "random_sequence.svh"
    `include "runall_sequence.svh"
    `include "mode_a_test.svh"
    `include "mode_b_test.svh"
    `include "random_test.svh"
    `include "runall_test.svh"
    


endpackage 