package alu_pkg;
    import uvm_pkg ::*;
    `include "uvm_macros.svh";
    `include "sequence_item.svh";
    `include "sequencer.svh";
    `include "driver.svh";
    `include "monitor.svh";
    `include "agent.svh";
    `include "base_sequence.svh";
    `include "reset_seq.svh";
    `include "mode_A_seq.svh";
    `include "mode_B_seq.svh";
    `include "scoreboard.svh";
    `include "coverage.svh";
    `include "env.svh";
    `include "base_test.svh";
    `include "mode_A_test.svh";
    `include "mode_B_test.svh";
    `include "full_test.svh";
    
endpackage 